module uop_fetch (
  input wire [128:0] insn,
  
);

endmodule 