module mem_read (
    
);
    
endmodule